////////////////////////////////////////////////////////////////////////////////////////////////////
// Filename:    problem6_cgrundey.v
// Author:      Colin Grundey
// Date:        13 March 2018
// Version:     1
// Description: Problem 6 solution

module problem6_cgrundey(parity_control, input_word, output_word);
  input parity_control; // 0 - odd, 1 - even
  input [7:0] input_word;
  output [8:0] output_word;


endmodule
